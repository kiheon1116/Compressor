class transaction;
  bit  [63:0] data [16];
  bit  valid;

endclass

