class transaction;
  bit  [63:0] data [16];
  bit  valid;
  bit  comp_flag;

endclass

